module top_module ( input a, input b, output out );
    mod_a mod1(a, b, out);
endmodule
